module Start ( input [4:0]	addr,
						output [63:0]	data
					 );

	parameter ADDR_WIDTH = 5;
   parameter DATA_WIDTH =  64;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:31][63:0] ROM = {
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000111110000000000000000000000000000000000,
64'b0000000000000000000000001101111000000000000000000000000000000000,
64'b0000000000000000000000011101111000000000000000000000000000000000,
64'b0000000000000000000000011111100000000000000000000000000000000000,
64'b0000000000000000000000011111000101010000000000000000000000000000,
64'b0000000000000000000000011111100000000000000000000000000000000000,
64'b0000000000000000000000011111111000000000000000000000000000000000,
64'b0000000000000000000000011111111000000000000000000000000000000000,
64'b0000000000000000000000001111110000000000000000000000000000000000,
64'b0000000000000000000000000011100000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000011100100010011111001110011100000000000000000000000000,
64'b0000000000010000110010000100001000010100000000000000000000000000,
64'b0000000000011000101010000100001100011100000000000000000000000000,
64'b0000000000010000100110000100001000011000000000000000000000000000,
64'b0000000000011100100010000100001110010100000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000
};

assign data = ROM[addr];

endmodule  
