module Sprites ( input [6:0]	addr,
						output [15:0]	data
					 );

	parameter ADDR_WIDTH = 7;
   parameter DATA_WIDTH =  16;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:95][DATA_WIDTH-1:0] ROM = {
		 16'b0000011111110000, // left x01
		 16'b0000111111111000,
		 16'b0001111111111100,
	    16'b0011111111111111,
		 16'b0011111111111110,
		 16'b0111111111111100,
		 16'b0111111111111000,
		 16'b0111111111100000,
		 16'b0111111111100000,
		 16'b0011111111111000,
		 16'b0011111111111100,
		 16'b0011111111111110,
		 16'b0011111111111111,
		 16'b0001111111111100,
		 16'b0000111111111000,
		 16'b0000011111110000,
		  
         
		16'b0000111111110000, // closed x02
		16'b0001111111111000,
		16'b0011111111111100,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0111111111111110,
		16'b0011111111111100,
		16'b0001111111111000,
		16'b0000111111110000,

		  16'b0000111111110000,
		  16'b0011111111111100,
		  16'b1110011111100111,
		  16'b1101101111011011,
		  16'b1110011111100111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111111111111111,
		  16'b1111001111100111,
		  16'b1110000111000011,
		  16'b1100000010000001,
		  
16'b0001000000001000, //up x04
16'b0001100000011000,
16'b0011110000111100,
16'b0111111001111110,
16'b1111111001111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b0111111111111110,
16'b0011111111111100,
16'b0001111111111000,
16'b0000000110000000,
16'b0000000000000000,

16'b0000000000000000, // down x05
16'b0000000110000000,
16'b0001111111111000,
16'b0011111111111100,
16'b0111111111111110,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111111111111,
16'b1111111001111111,
16'b0111111001111110,
16'b0011110000111100,
16'b0001100000011000,
16'b0001000000001000,

16'b0000111111100000, // right x06
16'b0001111111110000,
16'b0011111111111000,
16'b1111111111111100,
16'b0111111111111100,
16'b0011111111111110,
16'b0001111111111110,
16'b0000011111111110,
16'b0000011111111110,
16'b0001111111111110,
16'b0011111111111100,
16'b0111111111111100,
16'b1111111111111100,
16'b0011111111111000,
16'b0001111111110000,
16'b0000111111100000
        };

	assign data = ROM[addr];

endmodule  