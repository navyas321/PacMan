module Win ( input [4:0]	addr,
						output [63:0]	data
					 );

	parameter ADDR_WIDTH = 5;
   parameter DATA_WIDTH =  64;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:31][63:0] ROM = {
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000001111100000000000000000000000000000000000,
64'b0000000000000000000000001101111000000000000000000000000000000000,
64'b0000000000000000000000011101111000000000000000000000000000000000,
64'b0000000000000000000000011111100000000000000000000000000000000000,
64'b0000000000000000000000011111000000000000000000000000000000000000,
64'b0000000000000000000000011111100000000000000000000000000000000000,
64'b0000000000000000000000011111111000000000000000000000000000000000,
64'b0000000000000000000000011111111000000000000000000000000000000000,
64'b0000000000000000000000001111110000000000000000000000000000000000,
64'b0000000000000000000000000011100000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000010001001111001001000000010000010000010010010001000000000000,
64'b0000001010001001001001000000001000010000100010011001000000000000,
64'b0000000100001001001001000000000100101001000010010101000000000000,
64'b0000000100001001001001000000000011000101000010010011000000000000,
64'b0000000100001111001111000000000010000010000010010001000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000
};

assign data = ROM[addr];

endmodule  