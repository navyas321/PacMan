module End ( input [5:0]	addr,
						output [63:0]	data
					 );
parameter [0:31][63:0] ROM = {
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000100000000001000000000000000000000000000000,
64'b0000000000000000000000010111110010000000000000000000000000000000,
64'b0000000000000000000000001101111000000000000000000000000000000000,
64'b0000000000000000000000011101111000000000000000000000000000000000,
64'b0000000000000000000000011111100000000000000000000000000000000000,
64'b0000000000000000000000011111000000000000000000000000000000000000,
64'b0000000000000000000000011111100000000000000000000000000000000000,
64'b0000000000000000000000011111111000000000000000000000000000000000,
64'b0000000000000000000000011111111000000000000000000000000000000000,
64'b0000000000000000000000101111110100000000000000000000000000000000,
64'b0000000000000000000001000011100010000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000010001001111001001000000100000111100111100111110000000000000,
64'b0000001010001001001001000000100000100100100000100000000000000000,
64'b0000000100001001001001000000100000100100111100111110000000000000,
64'b0000000100001001001001000000100000100100000100100000000000000000,
64'b0000000100001111001111000000111100111100111100111110000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000,
64'b0000000000000000000000000000000000000000000000000000000000000000
};

assign data = ROM[addr];

endmodule  