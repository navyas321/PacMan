module testbench();

timeunit 10ns;	// Half clock cycle at 50 MHz
			// This is the amount of time represented by #1 
timeprecision 1ns;

// These signals are internal because the processor will be 
// instantiated as a submodule in testbench.
logic Clk = 0;
logic Reset;
logic [15:0]keyboard;
			//input logic pause
logic  pacDeath;
logic winsignal;
logic startscreen;
logic gamescreen;
			//output logic pausescreen,
logic gameoverscreen;
logic winscreen;

				
// A counter to count the instances where simulation results
// do no match with expected results


		
// Instantiating the DUT
// Make sure the module and signal names match with those in your design
FSM processor0(.*);	

// Toggle the clock
// #1 means wait for a delay of 1 timeunit
always begin : CLOCK_GENERATION
#1 Clk = ~Clk;
end

initial begin: CLOCK_INITIALIZATION
    Clk = 0;
end 

// Testing begins here
// The initial block is not synthesizable
// Everything happens sequentially inside an initial block
// as in a software program
initial begin: TEST_VECTORS
Reset = 0;		// Toggle Res
keyboard = 0;
pacDeath = 0;
winsignal = 0;

#2 Reset = 1;
#2 Reset = 0;
#2 keyboard = 8'h28;
#2 keyboard = 0;
#2 pacDeath = 1;
#2 pacDeath = 0;
#2 keyboard = 8'h2c;
#2 keyboard = 0;
#2 keyboard = 8'h28;
#2 keyboard = 0;
#2 winsignal = 1;
#2 winsignal = 0;
#2 keyboard = 8'h2c;
#2 keyboard = 0;

end
endmodule



